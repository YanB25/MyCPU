module REGISTER_FILE_TB(
);

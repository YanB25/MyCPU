`timescale 1ns/1ps

`include "head.v"
module REGISTER_FILE_TB(
);
    reg [DATA_WID - 1:0] data;
    initial begin
        


module REGEST_FILE (
);
    
